`define data_width 8
`define no_of_transactions 50
`define depth 16
